--************************************************************************************************
--  Generic AVR status register definitions.
--
--  Authors:
--      -- Kyle J. Temkin, Binghamton University, <ktemkin@binghamton.edu>
--************************************************************************************************

library ieee;
use ieee.std_logic_1164.all;

