--************************************************************************************************
--
-- AVR109-Compatible 
-- 
--
-- Authors include:
--     -Kyle J. Temkin, Binghamton University, <ktemkin@binghamton.edu>
--
--************************************************************************************************


library IEEE;
use IEEE.std_logic_1164.all;


entity avr109_programmer is

end avr109_programmer;

architecture Behavioral of avr109_programmer is

begin


end Behavioral;

